// Read only memory for spaceship RGB data storage

module shape_rom (clk, addr, data_out);
	input clk;
	input [7:0] addr;
	output reg [11:0] data_out;

	reg [11:0] rom [0:255];
	
	initial begin		// Fill rom with RGB values
		rom[0] = 12'h000;
		rom[1] = 12'h000;
		rom[2] = 12'h000;
		rom[3] = 12'h000;
		rom[4] = 12'h000;
		rom[5] = 12'h000;
		rom[6] = 12'h000;
		rom[7] = 12'h000;
		rom[8] = 12'h000;
		rom[9] = 12'h000;
		rom[10] = 12'h000;
		rom[11] = 12'h000;
		rom[12] = 12'h000;
		rom[13] = 12'h000;
		rom[14] = 12'h000;
		rom[15] = 12'h000;
		rom[16] = 12'h000;
		rom[17] = 12'h000;
		rom[18] = 12'hb2a;		// violet
		rom[19] = 12'haaa;		// silver
		rom[20] = 12'haaa;
		rom[21] = 12'haaa;
		rom[22] = 12'haaa;
		rom[23] = 12'hf80;		// orange
		rom[24] = 12'hf80;
		rom[25] = 12'h000;
		rom[26] = 12'h000;
		rom[27] = 12'h000;
		rom[28] = 12'h000;
		rom[29] = 12'h000;
		rom[30] = 12'h000;
		rom[31] = 12'h000;
		rom[32] = 12'h000;
		rom[33] = 12'h000;
		rom[34] = 12'h000;
		rom[35] = 12'hb2a;
		rom[36] = 12'h000;
		rom[37] = 12'h000;
		rom[38] = 12'h000;
		rom[39] = 12'h000;
		rom[40] = 12'h000;
		rom[41] = 12'h000;
		rom[42] = 12'h000;
		rom[43] = 12'h000;
		rom[44] = 12'h000;
		rom[45] = 12'h000;
		rom[46] = 12'h000;
		rom[47] = 12'h000;
		rom[48] = 12'hf80;
		rom[49] = 12'h333;	// dark gray
		rom[50] = 12'haaa;
		rom[51] = 12'haaa;
		rom[52] = 12'h000;
		rom[53] = 12'hb2a;
		rom[54] = 12'haaa;
		rom[55] = 12'haaa;
		rom[56] = 12'haaa;
		rom[57] = 12'hf80;
		rom[58] = 12'hf80;
		rom[59] = 12'h000;
		rom[60] = 12'h000;
		rom[61] = 12'h000;
		rom[62] = 12'h000;
		rom[63] = 12'h000;
		rom[64] = 12'hf80;
		rom[65] = 12'h333;
		rom[66] = 12'haaa;
		rom[67] = 12'haaa;
		rom[68] = 12'haaa;
		rom[69] = 12'haaa;
		rom[70] = 12'hb2a;
		rom[71] = 12'h000;
		rom[72] = 12'h000;
		rom[73] = 12'h000;
		rom[74] = 12'h000;
		rom[75] = 12'h000;
		rom[76] = 12'h000;
		rom[77] = 12'h000;
		rom[78] = 12'h000;
		rom[79] = 12'h000;
		rom[80] = 12'h000;
		rom[81] = 12'h000;
		rom[82] = 12'h000;
		rom[83] = 12'h000;
		rom[84] = 12'haaa;
		rom[85] = 12'haaa;
		rom[86] = 12'haaa;
		rom[87] = 12'haaa;
		rom[88] = 12'haaa;
		rom[89] = 12'h000;
		rom[90] = 12'h000;
		rom[91] = 12'h000;
		rom[92] = 12'h000;
		rom[93] = 12'h000;
		rom[94] = 12'h000;
		rom[95] = 12'h000;
		rom[96] = 12'h000;
		rom[97] = 12'h000;
		rom[98] = 12'h000;
		rom[99] = 12'haaa;
		rom[100] = 12'haaa;
		rom[101] = 12'h333;
		rom[102] = 12'h333;
		rom[103] = 12'haaa;
		rom[104] = 12'haaa;
		rom[105] = 12'haaa;
		rom[106] = 12'haaa;
		rom[107] = 12'haaa;
		rom[108] = 12'haaa;
		rom[109] = 12'haaa;
		rom[110] = 12'h000;
		rom[111] = 12'h000;
		rom[112] = 12'hf80;
		rom[113] = 12'h333;
		rom[114] = 12'haaa;
		rom[115] = 12'haaa;
		rom[116] = 12'haaa;
		rom[117] = 12'haaa;
		rom[118] = 12'h333;
		rom[119] = 12'h333;
		rom[120] = 12'haaa;
		rom[121] = 12'h333;
		rom[122] = 12'h333;
		rom[123] = 12'h333;
		rom[124] = 12'h333;
		rom[125] = 12'haaa;
		rom[126] = 12'haaa;
		rom[127] = 12'haaa;
		rom[128] = 12'hf80;
		rom[129] = 12'h333;
		rom[130] = 12'haaa;
		rom[131] = 12'haaa;
		rom[132] = 12'haaa;
		rom[133] = 12'haaa;
		rom[134] = 12'h333;
		rom[135] = 12'h333;
		rom[136] = 12'haaa;
		rom[137] = 12'h333;
		rom[138] = 12'h333;
		rom[139] = 12'h333;
		rom[140] = 12'h333;
		rom[141] = 12'haaa;
		rom[142] = 12'haaa;
		rom[143] = 12'haaa;
		rom[144] = 12'h000;
		rom[145] = 12'h000;
		rom[146] = 12'h000;
		rom[147] = 12'haaa;
		rom[148] = 12'haaa;
		rom[149] = 12'h333;
		rom[150] = 12'h333;
		rom[151] = 12'haaa;
		rom[152] = 12'haaa;
		rom[153] = 12'haaa;
		rom[154] = 12'haaa;
		rom[155] = 12'haaa;
		rom[156] = 12'haaa;
		rom[157] = 12'haaa;
		rom[158] = 12'h000;
		rom[159] = 12'h000;
		rom[160] = 12'h000;
		rom[161] = 12'h000;
		rom[162] = 12'h000;
		rom[163] = 12'h000;
		rom[164] = 12'haaa;
		rom[165] = 12'haaa;
		rom[166] = 12'haaa;
		rom[167] = 12'haaa;
		rom[168] = 12'haaa;
		rom[169] = 12'h000;
		rom[170] = 12'h000;
		rom[171] = 12'h000;
		rom[172] = 12'h000;
		rom[173] = 12'h000;
		rom[174] = 12'h000;
		rom[175] = 12'h000;
		rom[176] = 12'hf80;
		rom[177] = 12'h333;
		rom[178] = 12'haaa;
		rom[179] = 12'haaa;
		rom[180] = 12'haaa;
		rom[181] = 12'haaa;
		rom[182] = 12'hb2a;
		rom[183] = 12'h000;
		rom[184] = 12'h000;
		rom[185] = 12'h000;
		rom[186] = 12'h000;
		rom[187] = 12'h000;
		rom[188] = 12'h000;
		rom[189] = 12'h000;
		rom[190] = 12'h000;
		rom[191] = 12'h000;
		rom[192] = 12'hf80;
		rom[193] = 12'h333;
		rom[194] = 12'haaa;
		rom[195] = 12'haaa;
		rom[196] = 12'h000;
		rom[197] = 12'hb2a;
		rom[198] = 12'haaa;
		rom[199] = 12'haaa;
		rom[200] = 12'haaa;
		rom[201] = 12'hf80;
		rom[202] = 12'hf80;
		rom[203] = 12'h000;
		rom[204] = 12'h000;
		rom[205] = 12'h000;
		rom[206] = 12'h000;
		rom[207] = 12'h000;
		rom[208] = 12'h000;
		rom[209] = 12'h000;
		rom[210] = 12'h000;
		rom[211] = 12'hb2a;
		rom[212] = 12'h000;
		rom[213] = 12'h000;
		rom[214] = 12'h000;
		rom[215] = 12'h000;
		rom[216] = 12'h000;
		rom[217] = 12'h000;
		rom[218] = 12'h000;
		rom[219] = 12'h000;
		rom[220] = 12'h000;
		rom[221] = 12'h000;
		rom[222] = 12'h000;
		rom[223] = 12'h000;
		rom[224] = 12'h000;
		rom[225] = 12'h000;
		rom[226] = 12'hb2a;
		rom[227] = 12'haaa;
		rom[228] = 12'haaa;
		rom[229] = 12'haaa;
		rom[230] = 12'haaa;
		rom[231] = 12'hf80;
		rom[232] = 12'hf80;
		rom[233] = 12'h000;
		rom[234] = 12'h000;
		rom[235] = 12'h000;
		rom[236] = 12'h000;
		rom[237] = 12'h000;
		rom[238] = 12'h000;
		rom[239] = 12'h000;
		rom[240] = 12'h000;
		rom[241] = 12'h000;
		rom[242] = 12'h000;
		rom[243] = 12'h000;
		rom[244] = 12'h000;
		rom[245] = 12'h000;
		rom[246] = 12'h000;
		rom[247] = 12'h000;
		rom[248] = 12'h000;
		rom[249] = 12'h000;
		rom[250] = 12'h000;
		rom[251] = 12'h000;
		rom[252] = 12'h000;
		rom[253] = 12'h000;
		rom[254] = 12'h000;
		rom[255] = 12'h000;
	end				// Initial rom block
	
	always @ (posedge clk)			// Read rom every cycle
	begin
		data_out <= #1 rom[addr];
	end
endmodule